module cache_memory();

endmodule